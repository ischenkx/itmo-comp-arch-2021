module alu(srca, srcb, alucontrol, aluresult, zero);
  input [31:0] srca, srcb;
  input [2:0] alucontrol;
  output [31:0] aluresult;
  output zero;

  // TODO: implementation
endmodule
